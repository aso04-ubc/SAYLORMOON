module sha256(
    input logic clock,
    input logic reset,
    input logic start,
    input logic [511:0] block,
    output logic [255:0] digest,
    output logic finish
);

    function automatic logic [31:0] rotate_right(input logic[31:0] in, input int positions);
        // return {x[0], x[31:1]};
        return (in >> positions) | (in << (32-positions));
    endfunction

    function automatic logic [31:0] s0(input logic[31:0] in);
        return (rotate_right(in, 7) ^ rotate_right(in,18) ^ (in >> 3));
    endfunction

    function automatic logic [31:0] s1(input logic [31:0] in);
        return (rotate_right(in, 17) ^ rotate_right(in, 19) ^ (in >> 10));
    endfunction

    function automatic logic [31:0] choose(input logic [31:0] select, input logic [31:0] x, input logic [31:0] y);
        return (x & select) ^ (y & ~select);
    endfunction

    function automatic logic [31:0] majority (input logic [31:0] j, input logic [31:0] k, input logic [31:0] l);
        return (j & k) ^ (j & l) ^ (k & l);
    endfunction

    function automatic logic [31:0] S0 (input logic [31:0] in);
        return rotate_right(in, 2) ^ rotate_right(in, 13) ^ rotate_right(in, 22);
    endfunction

    function automatic logic [31:0] S1 (input logic [31:0] in);
        return rotate_right(in, 6) ^ rotate_right(in, 11) ^ rotate_right(in ,25);
    endfunction

    
    logic [31:0] temp1;
    logic [31:0] temp2;
    logic [31:0] W [0:63];

    logic [31:0] a, b, c, d, e, f, g, h;
    logic [31:0] H0, H1, H2, H3, H4, H5, H6, H7;
    logic [31:0] w_update;
    logic [6:0] timer;

    localparam logic [31:0] K [0:63] = '{
    32'h428a2f98, 32'h71374491, 32'hb5c0fbcf, 32'he9b5dba5, 32'h3956c25b, 32'h59f111f1, 32'h923f82a4, 32'hab1c5ed5,
    32'hd807aa98, 32'h12835b01, 32'h243185be, 32'h550c7dc3, 32'h72be5d74, 32'h80deb1fe, 32'h9bdc06a7, 32'hc19bf174,
    32'he49b69c1, 32'hefbe4786, 32'h0fc19dc6, 32'h240ca1cc, 32'h2de92c6f, 32'h4a7484aa, 32'h5cb0a9dc, 32'h76f988da,
    32'h983e5152, 32'ha831c66d, 32'hb00327c8, 32'hbf597fc7, 32'hc6e00bf3, 32'hd5a79147, 32'h06ca6351, 32'h14292967,
    32'h27b70a85, 32'h2e1b2138, 32'h4d2c6dfc, 32'h53380d13, 32'h650a7354, 32'h766a0abb, 32'h81c2c92e, 32'h92722c85,
    32'ha2bfe8a1, 32'ha81a664b, 32'hc24b8b70, 32'hc76c51a3, 32'hd192e819, 32'hd6990624, 32'hf40e3585, 32'h106aa070,
    32'h19a4c116, 32'h1e376c08, 32'h2748774c, 32'h34b0bcb5, 32'h391c0cb3, 32'h4ed8aa4a, 32'h5b9cca4f, 32'h682e6ff3,
    32'h748f82ee, 32'h78a5636f, 32'h84c87814, 32'h8cc70208, 32'h90befffa, 32'ha4506ceb, 32'hbef9a3f7, 32'hc67178f2
    };

    // anti pipeline hazard //
    assign temp1 = h + S1(e) + choose(e,f,g) + K[timer] + w_update;
    assign temp2 = S0(a) + majority(a,b,c);

    always_comb begin
        if (timer < 16) begin
            w_update = block[511 - timer * 32 -: 32];
        end else begin
            w_update = s1(W[timer-2]) + W[timer-7] + s0(W[timer-15]) + W[timer-16];
        end
    end
    // anti pipeline hazard //

    always_ff @(posedge clock or negedge reset) begin
        if (!reset) begin

            timer <= 7'd65;
            finish <= 0;

            H0 <= 32'h6a09e667;
            H1 <= 32'hbb67ae85;
            H2 <= 32'h3c6ef372;
            H3 <= 32'ha54ff53a;
            H4 <= 32'h510e527f;
            H5 <= 32'h9b05688c;
            H6 <= 32'h1f83d9ab;
            H7 <= 32'h5be0cd19;

        end else if (start && timer > 63) begin

            finish <= 0;
            timer <= 7'd0;

            a <= H0; b <= H1; c <= H2; d <= H3;
            e <= H4; f <= H5; g <= H6; h <= H7;

        end else if (timer < 64) begin

            W[timer] <= w_update;

            h <= g;
            g <= f;
            f <= e;
            e <= d + temp1;
            d <= c;
            c <= b;
            b <= a;
            a <= temp1 + temp2;

            timer <= timer + 1;

        end else if (timer == 64) begin

            H0 <= H0 + a; H1 <= H1 + b; H2 <= H2 + c; H3 <= H3 + d;
            H4 <= H4 + e; H5 <= H5 + f; H6 <= H6 + g; H7 <= H7 + h;

            finish <= 1;
            timer <= 7'd65;
        
        end
    end

    assign digest = {H0, H1, H2, H3, H4, H5, H6, H7};

endmodule